module brick_logic(
	input [9:0] col_x1, col_x2, col_y1, col_y2,
	
	input collided_1, collided_2
	);
