module loadFSM(
	input resetn,
	input clk,
	input [9:0]selection,
	
	output 
	);